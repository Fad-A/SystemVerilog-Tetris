// ## Fadi Ajaj ## 


Module replaceRow(input logic[19:0] inputRow, output logic[19:0] outputRow)

endmodule